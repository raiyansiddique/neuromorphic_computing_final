magic
tech sky130A
timestamp 1702611732
<< nwell >>
rect -125 -65 2255 275
<< nmos >>
rect -55 -560 -5 -260
rect 45 -560 95 -260
rect 225 -560 275 -260
rect 325 -560 375 -260
rect 425 -560 475 -260
rect 525 -560 575 -260
rect 625 -560 675 -260
rect 805 -560 855 -260
rect 1055 -560 1105 -260
rect 1235 -560 1285 -260
rect 1335 -560 1385 -260
rect 1435 -560 1485 -260
rect 1535 -560 1585 -260
rect 1635 -560 1685 -260
rect 1735 -560 1785 -260
rect 1835 -560 1885 -260
rect 1935 -560 1985 -260
rect 2035 -560 2085 -260
rect 2135 -560 2185 -260
<< pmos >>
rect -55 -45 -5 255
rect 45 -45 95 255
rect 145 -45 195 255
rect 245 -45 295 255
rect 345 -45 395 255
rect 445 -45 495 255
rect 545 -45 595 255
rect 645 -45 695 255
rect 745 -45 795 255
rect 845 -45 895 255
rect 1075 -45 1125 255
rect 1275 -45 1325 255
rect 1455 -45 1505 255
rect 1555 -45 1605 255
rect 1735 -45 1785 255
rect 1835 -45 1885 255
rect 1935 -45 1985 255
rect 2035 -45 2085 255
rect 2135 -45 2185 255
<< ndiff >>
rect -105 -275 -55 -260
rect -105 -545 -90 -275
rect -70 -545 -55 -275
rect -105 -560 -55 -545
rect -5 -275 45 -260
rect -5 -545 10 -275
rect 30 -545 45 -275
rect -5 -560 45 -545
rect 95 -275 145 -260
rect 95 -545 110 -275
rect 130 -545 145 -275
rect 95 -560 145 -545
rect 175 -275 225 -260
rect 175 -545 190 -275
rect 210 -545 225 -275
rect 175 -560 225 -545
rect 275 -275 325 -260
rect 275 -545 290 -275
rect 310 -545 325 -275
rect 275 -560 325 -545
rect 375 -275 425 -260
rect 375 -545 390 -275
rect 410 -545 425 -275
rect 375 -560 425 -545
rect 475 -275 525 -260
rect 475 -545 490 -275
rect 510 -545 525 -275
rect 475 -560 525 -545
rect 575 -275 625 -260
rect 575 -545 590 -275
rect 610 -545 625 -275
rect 575 -560 625 -545
rect 675 -275 725 -260
rect 675 -545 690 -275
rect 710 -545 725 -275
rect 675 -560 725 -545
rect 755 -275 805 -260
rect 755 -545 770 -275
rect 790 -545 805 -275
rect 755 -560 805 -545
rect 855 -275 905 -260
rect 855 -545 870 -275
rect 890 -545 905 -275
rect 855 -560 905 -545
rect 1005 -275 1055 -260
rect 1005 -545 1020 -275
rect 1040 -545 1055 -275
rect 1005 -560 1055 -545
rect 1105 -275 1155 -260
rect 1105 -545 1120 -275
rect 1140 -545 1155 -275
rect 1105 -560 1155 -545
rect 1185 -275 1235 -260
rect 1185 -545 1200 -275
rect 1220 -545 1235 -275
rect 1185 -560 1235 -545
rect 1285 -275 1335 -260
rect 1285 -545 1300 -275
rect 1320 -545 1335 -275
rect 1285 -560 1335 -545
rect 1385 -275 1435 -260
rect 1385 -545 1400 -275
rect 1420 -545 1435 -275
rect 1385 -560 1435 -545
rect 1485 -275 1535 -260
rect 1485 -545 1500 -275
rect 1520 -545 1535 -275
rect 1485 -560 1535 -545
rect 1585 -275 1635 -260
rect 1585 -545 1600 -275
rect 1620 -545 1635 -275
rect 1585 -560 1635 -545
rect 1685 -275 1735 -260
rect 1685 -545 1700 -275
rect 1720 -545 1735 -275
rect 1685 -560 1735 -545
rect 1785 -275 1835 -260
rect 1785 -545 1800 -275
rect 1820 -545 1835 -275
rect 1785 -560 1835 -545
rect 1885 -275 1935 -260
rect 1885 -545 1900 -275
rect 1920 -545 1935 -275
rect 1885 -560 1935 -545
rect 1985 -275 2035 -260
rect 1985 -545 2000 -275
rect 2020 -545 2035 -275
rect 1985 -560 2035 -545
rect 2085 -275 2135 -260
rect 2085 -545 2100 -275
rect 2120 -545 2135 -275
rect 2085 -560 2135 -545
rect 2185 -275 2235 -260
rect 2185 -545 2200 -275
rect 2220 -545 2235 -275
rect 2185 -560 2235 -545
<< pdiff >>
rect -105 240 -55 255
rect -105 -30 -90 240
rect -70 -30 -55 240
rect -105 -45 -55 -30
rect -5 240 45 255
rect -5 -30 10 240
rect 30 -30 45 240
rect -5 -45 45 -30
rect 95 240 145 255
rect 95 -30 110 240
rect 130 -30 145 240
rect 95 -45 145 -30
rect 195 240 245 255
rect 195 -30 210 240
rect 230 -30 245 240
rect 195 -45 245 -30
rect 295 240 345 255
rect 295 -30 310 240
rect 330 -30 345 240
rect 295 -45 345 -30
rect 395 240 445 255
rect 395 -30 410 240
rect 430 -30 445 240
rect 395 -45 445 -30
rect 495 240 545 255
rect 495 -30 510 240
rect 530 -30 545 240
rect 495 -45 545 -30
rect 595 240 645 255
rect 595 -30 610 240
rect 630 -30 645 240
rect 595 -45 645 -30
rect 695 240 745 255
rect 695 -30 710 240
rect 730 -30 745 240
rect 695 -45 745 -30
rect 795 240 845 255
rect 795 -30 810 240
rect 830 -30 845 240
rect 795 -45 845 -30
rect 895 240 945 255
rect 895 -30 910 240
rect 930 -30 945 240
rect 895 -45 945 -30
rect 1025 240 1075 255
rect 1025 -30 1040 240
rect 1060 -30 1075 240
rect 1025 -45 1075 -30
rect 1125 240 1175 255
rect 1125 -30 1140 240
rect 1160 -30 1175 240
rect 1125 -45 1175 -30
rect 1225 240 1275 255
rect 1225 -30 1240 240
rect 1260 -30 1275 240
rect 1225 -45 1275 -30
rect 1325 240 1375 255
rect 1325 -30 1340 240
rect 1360 -30 1375 240
rect 1325 -45 1375 -30
rect 1405 240 1455 255
rect 1405 -30 1420 240
rect 1440 -30 1455 240
rect 1405 -45 1455 -30
rect 1505 240 1555 255
rect 1505 -30 1520 240
rect 1540 -30 1555 240
rect 1505 -45 1555 -30
rect 1605 240 1655 255
rect 1605 -30 1620 240
rect 1640 -30 1655 240
rect 1605 -45 1655 -30
rect 1685 240 1735 255
rect 1685 -30 1700 240
rect 1720 -30 1735 240
rect 1685 -45 1735 -30
rect 1785 240 1835 255
rect 1785 -30 1800 240
rect 1820 -30 1835 240
rect 1785 -45 1835 -30
rect 1885 240 1935 255
rect 1885 -30 1900 240
rect 1920 -30 1935 240
rect 1885 -45 1935 -30
rect 1985 240 2035 255
rect 1985 -30 2000 240
rect 2020 -30 2035 240
rect 1985 -45 2035 -30
rect 2085 240 2135 255
rect 2085 -30 2100 240
rect 2120 -30 2135 240
rect 2085 -45 2135 -30
rect 2185 240 2235 255
rect 2185 -30 2200 240
rect 2220 -30 2235 240
rect 2185 -45 2235 -30
<< ndiffc >>
rect -90 -545 -70 -275
rect 10 -545 30 -275
rect 110 -545 130 -275
rect 190 -545 210 -275
rect 290 -545 310 -275
rect 390 -545 410 -275
rect 490 -545 510 -275
rect 590 -545 610 -275
rect 690 -545 710 -275
rect 770 -545 790 -275
rect 870 -545 890 -275
rect 1020 -545 1040 -275
rect 1120 -545 1140 -275
rect 1200 -545 1220 -275
rect 1300 -545 1320 -275
rect 1400 -545 1420 -275
rect 1500 -545 1520 -275
rect 1600 -545 1620 -275
rect 1700 -545 1720 -275
rect 1800 -545 1820 -275
rect 1900 -545 1920 -275
rect 2000 -545 2020 -275
rect 2100 -545 2120 -275
rect 2200 -545 2220 -275
<< pdiffc >>
rect -90 -30 -70 240
rect 10 -30 30 240
rect 110 -30 130 240
rect 210 -30 230 240
rect 310 -30 330 240
rect 410 -30 430 240
rect 510 -30 530 240
rect 610 -30 630 240
rect 710 -30 730 240
rect 810 -30 830 240
rect 910 -30 930 240
rect 1040 -30 1060 240
rect 1140 -30 1160 240
rect 1240 -30 1260 240
rect 1340 -30 1360 240
rect 1420 -30 1440 240
rect 1520 -30 1540 240
rect 1620 -30 1640 240
rect 1700 -30 1720 240
rect 1800 -30 1820 240
rect 1900 -30 1920 240
rect 2000 -30 2020 240
rect 2100 -30 2120 240
rect 2200 -30 2220 240
<< psubdiff >>
rect 955 -275 1005 -260
rect 955 -545 970 -275
rect 990 -545 1005 -275
rect 955 -560 1005 -545
<< nsubdiff >>
rect 975 240 1025 255
rect 975 -30 990 240
rect 1010 -30 1025 240
rect 975 -45 1025 -30
<< psubdiffcont >>
rect 970 -545 990 -275
<< nsubdiffcont >>
rect 990 -30 1010 240
<< poly >>
rect 155 300 195 310
rect 155 280 165 300
rect 185 280 195 300
rect 155 270 195 280
rect 255 300 295 310
rect 255 280 265 300
rect 285 280 295 300
rect 255 270 295 280
rect 355 300 395 310
rect 355 280 365 300
rect 385 280 395 300
rect 355 270 395 280
rect -55 255 -5 270
rect 45 255 95 270
rect 145 255 195 270
rect 245 255 295 270
rect 345 255 395 270
rect 445 300 485 310
rect 445 280 455 300
rect 475 280 485 300
rect 445 270 485 280
rect 545 300 585 310
rect 545 280 555 300
rect 575 280 585 300
rect 545 270 585 280
rect 645 300 685 310
rect 645 280 655 300
rect 675 280 685 300
rect 645 270 685 280
rect 1075 300 1115 310
rect 1075 280 1085 300
rect 1105 280 1115 300
rect 1075 270 1115 280
rect 1275 300 1315 310
rect 1275 280 1285 300
rect 1305 280 1315 300
rect 1275 270 1315 280
rect 1410 300 1450 310
rect 1410 280 1420 300
rect 1440 285 1450 300
rect 2190 300 2230 310
rect 2190 285 2200 300
rect 1440 280 1605 285
rect 1410 270 1605 280
rect 445 255 495 270
rect 545 255 595 270
rect 645 255 695 270
rect 745 255 795 270
rect 845 255 895 270
rect 1075 255 1125 270
rect 1275 255 1325 270
rect 1455 255 1505 270
rect 1555 255 1605 270
rect 1735 280 2200 285
rect 2220 280 2230 300
rect 1735 270 2230 280
rect 1735 255 1785 270
rect 1835 255 1885 270
rect 1935 255 1985 270
rect 2035 255 2085 270
rect 2135 255 2185 270
rect -55 -60 -5 -45
rect 45 -60 95 -45
rect 145 -60 195 -45
rect 245 -60 295 -45
rect -55 -75 95 -60
rect 80 -85 95 -75
rect 345 -85 395 -45
rect 445 -85 495 -45
rect 545 -60 595 -45
rect 645 -60 695 -45
rect 745 -60 795 -45
rect 845 -60 895 -45
rect 1075 -60 1125 -45
rect 1275 -60 1325 -45
rect 1455 -60 1505 -45
rect 1555 -60 1605 -45
rect 1735 -60 1785 -45
rect 1835 -60 1885 -45
rect 1935 -60 1985 -45
rect 2035 -60 2085 -45
rect 2135 -60 2185 -45
rect 745 -75 895 -60
rect 920 -75 1095 -60
rect 745 -85 760 -75
rect 80 -100 760 -85
rect 620 -165 660 -155
rect 620 -185 630 -165
rect 650 -180 660 -165
rect 820 -165 860 -155
rect 820 -180 830 -165
rect 650 -185 830 -180
rect 850 -185 860 -165
rect 620 -195 860 -185
rect 920 -230 940 -75
rect 990 -110 1030 -100
rect 990 -130 1000 -110
rect 1020 -125 1030 -110
rect 1090 -110 1130 -100
rect 1090 -125 1100 -110
rect 1020 -130 1100 -125
rect 1120 -130 1130 -110
rect 990 -140 1130 -130
rect 1440 -110 1580 -100
rect 1440 -130 1450 -110
rect 1470 -115 1550 -110
rect 1470 -130 1480 -115
rect 1440 -140 1480 -130
rect 1540 -130 1550 -115
rect 1570 -130 1580 -110
rect 1540 -140 1580 -130
rect 990 -175 1140 -165
rect 990 -195 1000 -175
rect 1020 -180 1110 -175
rect 1020 -195 1030 -180
rect 990 -205 1030 -195
rect 1100 -195 1110 -180
rect 1130 -195 1140 -175
rect 1100 -205 1140 -195
rect 1370 -220 2050 -205
rect 1370 -230 1385 -220
rect 805 -245 1105 -230
rect -55 -260 -5 -245
rect 45 -260 95 -245
rect 225 -260 275 -245
rect 325 -260 375 -245
rect 425 -260 475 -245
rect 525 -260 575 -245
rect 625 -260 675 -245
rect 805 -260 855 -245
rect 1055 -260 1105 -245
rect 1235 -245 1385 -230
rect 1235 -260 1285 -245
rect 1335 -260 1385 -245
rect 1435 -260 1485 -245
rect 1535 -260 1585 -245
rect 1635 -260 1685 -220
rect 1735 -260 1785 -220
rect 2035 -230 2050 -220
rect 2035 -245 2185 -230
rect 1835 -260 1885 -245
rect 1935 -260 1985 -245
rect 2035 -260 2085 -245
rect 2135 -260 2185 -245
rect -55 -575 -5 -560
rect 45 -575 95 -560
rect -100 -585 95 -575
rect -100 -605 -90 -585
rect -70 -590 95 -585
rect 225 -575 275 -560
rect 325 -575 375 -560
rect 425 -575 475 -560
rect 525 -575 575 -560
rect 625 -575 675 -560
rect 805 -575 855 -560
rect 1055 -575 1105 -560
rect 1235 -575 1285 -560
rect 1335 -575 1385 -560
rect 1435 -575 1485 -560
rect 1535 -575 1585 -560
rect 1635 -575 1685 -560
rect 225 -585 720 -575
rect 225 -590 690 -585
rect -70 -605 -60 -590
rect -100 -615 -60 -605
rect 680 -605 690 -590
rect 710 -605 720 -585
rect 680 -615 720 -605
rect 1445 -585 1485 -575
rect 1445 -605 1455 -585
rect 1475 -605 1485 -585
rect 1445 -615 1485 -605
rect 1545 -585 1585 -575
rect 1545 -605 1555 -585
rect 1575 -605 1585 -585
rect 1545 -615 1585 -605
rect 1645 -585 1685 -575
rect 1645 -605 1655 -585
rect 1675 -605 1685 -585
rect 1645 -615 1685 -605
rect 1735 -575 1785 -560
rect 1835 -575 1885 -560
rect 1935 -575 1985 -560
rect 2035 -575 2085 -560
rect 2135 -575 2185 -560
rect 1735 -585 1775 -575
rect 1735 -605 1745 -585
rect 1765 -605 1775 -585
rect 1735 -615 1775 -605
rect 1835 -585 1875 -575
rect 1835 -605 1845 -585
rect 1865 -605 1875 -585
rect 1835 -615 1875 -605
rect 1935 -585 1975 -575
rect 1935 -605 1945 -585
rect 1965 -605 1975 -585
rect 1935 -615 1975 -605
<< polycont >>
rect 165 280 185 300
rect 265 280 285 300
rect 365 280 385 300
rect 455 280 475 300
rect 555 280 575 300
rect 655 280 675 300
rect 1085 280 1105 300
rect 1285 280 1305 300
rect 1420 280 1440 300
rect 2200 280 2220 300
rect 630 -185 650 -165
rect 830 -185 850 -165
rect 1000 -130 1020 -110
rect 1100 -130 1120 -110
rect 1450 -130 1470 -110
rect 1550 -130 1570 -110
rect 1000 -195 1020 -175
rect 1110 -195 1130 -175
rect -90 -605 -70 -585
rect 690 -605 710 -585
rect 1455 -605 1475 -585
rect 1555 -605 1575 -585
rect 1655 -605 1675 -585
rect 1745 -605 1765 -585
rect 1845 -605 1865 -585
rect 1945 -605 1965 -585
<< locali >>
rect 155 300 195 310
rect 155 280 165 300
rect 185 280 195 300
rect 155 270 195 280
rect 255 300 295 310
rect 255 280 265 300
rect 285 280 295 300
rect 255 270 295 280
rect 355 300 485 310
rect 355 280 365 300
rect 385 290 455 300
rect 385 280 395 290
rect 355 270 395 280
rect 445 280 455 290
rect 475 280 485 300
rect 445 270 485 280
rect 545 300 585 310
rect 545 280 555 300
rect 575 280 585 300
rect 545 270 585 280
rect 645 300 685 310
rect 645 280 655 300
rect 675 280 685 300
rect 645 270 685 280
rect 1075 300 1115 310
rect 1075 280 1085 300
rect 1105 280 1115 300
rect 1275 300 1315 310
rect 1275 290 1285 300
rect 1075 270 1115 280
rect 1150 280 1285 290
rect 1305 280 1315 300
rect 1150 270 1315 280
rect 1410 300 1450 310
rect 1410 280 1420 300
rect 1440 280 1450 300
rect 1410 270 1450 280
rect 2190 300 2230 310
rect 2190 280 2200 300
rect 2220 280 2230 300
rect 2190 270 2230 280
rect 1150 250 1170 270
rect 1410 250 1430 270
rect 2210 250 2230 270
rect -100 240 -60 250
rect -100 -30 -90 240
rect -70 -30 -60 240
rect -100 -40 -60 -30
rect 0 240 40 250
rect 0 -30 10 240
rect 30 -30 40 240
rect 0 -40 40 -30
rect 100 240 140 250
rect 100 -30 110 240
rect 130 -30 140 240
rect 100 -40 140 -30
rect 200 240 240 250
rect 200 -30 210 240
rect 230 -30 240 240
rect 200 -40 240 -30
rect 300 240 340 250
rect 300 -30 310 240
rect 330 -30 340 240
rect 300 -40 340 -30
rect 400 240 440 250
rect 400 -30 410 240
rect 430 -30 440 240
rect 400 -40 440 -30
rect 500 240 540 250
rect 500 -30 510 240
rect 530 -30 540 240
rect 500 -40 540 -30
rect 600 240 640 250
rect 600 -30 610 240
rect 630 -30 640 240
rect 600 -40 640 -30
rect 700 240 740 250
rect 700 -30 710 240
rect 730 -30 740 240
rect 700 -40 740 -30
rect 800 240 840 250
rect 800 -30 810 240
rect 830 -30 840 240
rect 800 -40 840 -30
rect 900 240 940 250
rect 900 -30 910 240
rect 930 -30 940 240
rect 900 -40 940 -30
rect 980 240 1070 250
rect 980 -30 990 240
rect 1010 -30 1040 240
rect 1060 -30 1070 240
rect 980 -40 1070 -30
rect 1130 240 1170 250
rect 1130 -30 1140 240
rect 1160 -30 1170 240
rect 1130 -40 1170 -30
rect 1230 240 1270 250
rect 1230 -30 1240 240
rect 1260 -30 1270 240
rect 1230 -40 1270 -30
rect 1330 240 1370 250
rect 1330 -30 1340 240
rect 1360 -30 1370 240
rect 1330 -40 1370 -30
rect 1410 240 1450 250
rect 1410 -30 1420 240
rect 1440 -30 1450 240
rect 1410 -40 1450 -30
rect 1510 240 1550 250
rect 1510 -30 1520 240
rect 1540 -30 1550 240
rect 1510 -40 1550 -30
rect 1610 240 1650 250
rect 1610 -30 1620 240
rect 1640 -30 1650 240
rect 1610 -40 1650 -30
rect 1690 240 1730 250
rect 1690 -30 1700 240
rect 1720 -30 1730 240
rect 1690 -40 1730 -30
rect 1790 240 1830 250
rect 1790 -30 1800 240
rect 1820 -30 1830 240
rect 1790 -40 1830 -30
rect 1890 240 1930 250
rect 1890 -30 1900 240
rect 1920 -30 1930 240
rect 1890 -40 1930 -30
rect 1990 240 2030 250
rect 1990 -30 2000 240
rect 2020 -30 2030 240
rect 1990 -40 2030 -30
rect 2090 240 2130 250
rect 2090 -30 2100 240
rect 2120 -30 2130 240
rect 2090 -40 2130 -30
rect 2190 240 2230 250
rect 2190 -30 2200 240
rect 2220 -30 2230 240
rect 2190 -40 2230 -30
rect -80 -75 -60 -40
rect 120 -75 140 -40
rect -80 -95 140 -75
rect 210 -115 230 -40
rect -80 -135 230 -115
rect 610 -115 630 -40
rect 700 -75 720 -40
rect 900 -75 920 -40
rect 1130 -60 1150 -40
rect 700 -95 920 -75
rect 1050 -80 1150 -60
rect 990 -110 1030 -100
rect 990 -115 1000 -110
rect 610 -135 700 -115
rect -80 -265 -60 -135
rect 620 -165 660 -155
rect 620 -175 630 -165
rect 480 -185 630 -175
rect 650 -185 660 -165
rect 480 -195 660 -185
rect 480 -225 500 -195
rect 120 -245 500 -225
rect 120 -265 140 -245
rect 280 -265 300 -245
rect 480 -265 500 -245
rect 680 -265 700 -135
rect 780 -130 1000 -115
rect 1020 -130 1030 -110
rect 780 -135 1030 -130
rect 780 -265 800 -135
rect 990 -140 1030 -135
rect 820 -165 860 -155
rect 820 -185 830 -165
rect 850 -175 860 -165
rect 990 -175 1030 -165
rect 850 -185 1000 -175
rect 820 -195 1000 -185
rect 1020 -195 1030 -175
rect -100 -275 -60 -265
rect -100 -545 -90 -275
rect -70 -545 -60 -275
rect -100 -555 -60 -545
rect 0 -275 40 -265
rect 0 -545 10 -275
rect 30 -545 40 -275
rect 0 -555 40 -545
rect 100 -275 140 -265
rect 100 -545 110 -275
rect 130 -545 140 -275
rect 100 -555 140 -545
rect 180 -275 220 -265
rect 180 -545 190 -275
rect 210 -545 220 -275
rect 180 -555 220 -545
rect 280 -275 320 -265
rect 280 -545 290 -275
rect 310 -545 320 -275
rect 280 -555 320 -545
rect 380 -275 420 -265
rect 380 -545 390 -275
rect 410 -545 420 -275
rect 380 -555 420 -545
rect 480 -275 520 -265
rect 480 -545 490 -275
rect 510 -545 520 -275
rect 480 -555 520 -545
rect 580 -275 620 -265
rect 580 -545 590 -275
rect 610 -545 620 -275
rect 580 -555 620 -545
rect 680 -275 720 -265
rect 680 -545 690 -275
rect 710 -545 720 -275
rect 680 -555 720 -545
rect 760 -275 800 -265
rect 760 -545 770 -275
rect 790 -545 800 -275
rect 760 -555 800 -545
rect 860 -265 880 -195
rect 990 -205 1030 -195
rect 1050 -225 1070 -80
rect 1230 -100 1250 -40
rect 1090 -110 1250 -100
rect 1090 -130 1100 -110
rect 1120 -120 1250 -110
rect 1330 -100 1350 -40
rect 1410 -60 1430 -40
rect 1630 -60 1650 -40
rect 1790 -60 1810 -40
rect 1990 -60 2010 -40
rect 1410 -80 1520 -60
rect 1330 -110 1480 -100
rect 1330 -120 1450 -110
rect 1120 -130 1130 -120
rect 1090 -140 1130 -130
rect 1330 -140 1350 -120
rect 1440 -130 1450 -120
rect 1470 -130 1480 -110
rect 1440 -140 1480 -130
rect 1150 -160 1350 -140
rect 1150 -165 1170 -160
rect 1100 -175 1170 -165
rect 1100 -195 1110 -175
rect 1130 -185 1170 -175
rect 1130 -195 1140 -185
rect 1100 -205 1140 -195
rect 1050 -245 1130 -225
rect 1110 -265 1130 -245
rect 1210 -230 1430 -210
rect 1210 -265 1230 -230
rect 1410 -265 1430 -230
rect 1500 -265 1520 -80
rect 1630 -80 2010 -60
rect 1630 -100 1650 -80
rect 2190 -100 2210 -40
rect 1540 -110 1650 -100
rect 1540 -130 1550 -110
rect 1570 -120 1650 -110
rect 1900 -120 2210 -100
rect 1570 -130 1580 -120
rect 1540 -140 1580 -130
rect 1900 -265 1920 -120
rect 1990 -230 2210 -210
rect 1990 -265 2010 -230
rect 2190 -265 2210 -230
rect 860 -275 900 -265
rect 860 -545 870 -275
rect 890 -545 900 -275
rect 860 -555 900 -545
rect 960 -275 1050 -265
rect 960 -545 970 -275
rect 990 -545 1020 -275
rect 1040 -545 1050 -275
rect 960 -555 1050 -545
rect 1110 -275 1150 -265
rect 1110 -545 1120 -275
rect 1140 -545 1150 -275
rect 1110 -555 1150 -545
rect 1190 -275 1230 -265
rect 1190 -545 1200 -275
rect 1220 -545 1230 -275
rect 1190 -555 1230 -545
rect 1290 -275 1330 -265
rect 1290 -545 1300 -275
rect 1320 -545 1330 -275
rect 1290 -555 1330 -545
rect 1390 -275 1430 -265
rect 1390 -545 1400 -275
rect 1420 -545 1430 -275
rect 1390 -555 1430 -545
rect 1490 -275 1530 -265
rect 1490 -545 1500 -275
rect 1520 -545 1530 -275
rect 1490 -555 1530 -545
rect 1590 -275 1630 -265
rect 1590 -545 1600 -275
rect 1620 -545 1630 -275
rect 1590 -555 1630 -545
rect 1690 -275 1730 -265
rect 1690 -545 1700 -275
rect 1720 -545 1730 -275
rect 1690 -555 1730 -545
rect 1790 -275 1830 -265
rect 1790 -545 1800 -275
rect 1820 -545 1830 -275
rect 1790 -555 1830 -545
rect 1890 -275 1930 -265
rect 1890 -545 1900 -275
rect 1920 -545 1930 -275
rect 1890 -555 1930 -545
rect 1990 -275 2030 -265
rect 1990 -545 2000 -275
rect 2020 -545 2030 -275
rect 1990 -555 2030 -545
rect 2090 -275 2130 -265
rect 2090 -545 2100 -275
rect 2120 -545 2130 -275
rect 2090 -555 2130 -545
rect 2190 -275 2230 -265
rect 2190 -545 2200 -275
rect 2220 -545 2230 -275
rect 2190 -555 2230 -545
rect -100 -575 -80 -555
rect 700 -575 720 -555
rect -100 -585 -60 -575
rect -100 -605 -90 -585
rect -70 -605 -60 -585
rect -100 -615 -60 -605
rect 680 -585 720 -575
rect 680 -605 690 -585
rect 710 -605 720 -585
rect 680 -615 720 -605
rect 780 -615 800 -555
rect 1445 -585 1485 -575
rect 1445 -605 1455 -585
rect 1475 -605 1485 -585
rect 1445 -615 1485 -605
rect 1545 -585 1585 -575
rect 1545 -605 1555 -585
rect 1575 -605 1585 -585
rect 1545 -615 1585 -605
rect 1645 -585 1685 -575
rect 1645 -605 1655 -585
rect 1675 -595 1685 -585
rect 1735 -585 1775 -575
rect 1735 -595 1745 -585
rect 1675 -605 1745 -595
rect 1765 -605 1775 -585
rect 1645 -615 1775 -605
rect 1835 -585 1875 -575
rect 1835 -605 1845 -585
rect 1865 -605 1875 -585
rect 1835 -615 1875 -605
rect 1935 -585 1975 -575
rect 1935 -605 1945 -585
rect 1965 -605 1975 -585
rect 1935 -615 1975 -605
<< viali >>
rect 10 -30 30 240
rect 410 -30 430 240
rect 810 -30 830 240
rect 990 -30 1010 240
rect 1040 -30 1060 240
rect 1520 -30 1540 240
rect 1700 -30 1720 240
rect 1900 -30 1920 240
rect 2100 -30 2120 240
rect 10 -545 30 -275
rect 190 -545 210 -275
rect 390 -545 410 -275
rect 590 -545 610 -275
rect 970 -545 990 -275
rect 1020 -545 1040 -275
rect 1300 -545 1320 -275
rect 1700 -545 1720 -275
rect 2100 -545 2120 -275
<< metal1 >>
rect -105 240 2235 255
rect -105 -30 10 240
rect 30 -30 410 240
rect 430 -30 810 240
rect 830 -30 990 240
rect 1010 -30 1040 240
rect 1060 -30 1520 240
rect 1540 -30 1700 240
rect 1720 -30 1900 240
rect 1920 -30 2100 240
rect 2120 -30 2235 240
rect -105 -45 2235 -30
rect -105 -275 2235 -260
rect -105 -545 10 -275
rect 30 -545 190 -275
rect 210 -545 390 -275
rect 410 -545 590 -275
rect 610 -545 970 -275
rect 990 -545 1020 -275
rect 1040 -545 1300 -275
rect 1320 -545 1700 -275
rect 1720 -545 2100 -275
rect 2120 -545 2235 -275
rect -105 -560 2235 -545
<< labels >>
rlabel locali 175 310 175 310 1 W1m
port 1 n
rlabel locali 275 310 275 310 1 W0m
port 2 n
rlabel locali 565 310 565 310 1 W2m
port 4 n
rlabel locali 665 310 665 310 1 W3m
port 5 n
rlabel locali 1465 -615 1465 -615 5 W1p
port 10 s
rlabel locali 1565 -615 1565 -615 5 W0p
port 11 s
rlabel locali 1855 -615 1855 -615 5 W2p
port 13 s
rlabel locali 1955 -615 1955 -615 5 W3p
port 14 s
rlabel metal1 -105 105 -105 105 7 VP
port 6 w
rlabel locali 420 310 420 310 1 VBP
port 3 n
rlabel locali 1710 -615 1710 -615 5 VBN
port 12 s
rlabel locali 790 -615 790 -615 5 IOUT
port 8 s
rlabel metal1 -105 -410 -105 -410 7 VN
port 15 w
rlabel locali 1095 310 1095 310 1 SPKIN
port 9 s
<< end >>
