magic
tech sky130A
timestamp 1702443510
<< nwell >>
rect -27 2513 1035 2641
rect -28 2474 1035 2513
rect -28 2177 308 2474
rect 89 2036 307 2177
rect 554 2034 1790 2274
<< nmos >>
rect 710 2360 1310 2390
rect 1375 2360 1825 2375
rect 425 2170 440 2270
rect 1876 2079 2076 2379
rect 0 0 2000 2000
<< pmos >>
rect 371 2542 971 2572
rect -10 2245 290 2445
rect 159 2054 174 2154
rect 572 2104 1772 2154
<< ndiff >>
rect 710 2428 1310 2440
rect 710 2403 724 2428
rect 1293 2403 1310 2428
rect 710 2390 1310 2403
rect 1375 2413 1825 2425
rect 1375 2389 1395 2413
rect 1807 2389 1825 2413
rect 1375 2375 1825 2389
rect 1876 2419 2076 2429
rect 1876 2393 1890 2419
rect 2061 2393 2076 2419
rect 1876 2379 2076 2393
rect 710 2348 1310 2360
rect 710 2323 723 2348
rect 1292 2323 1310 2348
rect 710 2310 1310 2323
rect 1375 2347 1825 2360
rect 1375 2323 1395 2347
rect 1807 2323 1825 2347
rect 1375 2310 1825 2323
rect 375 2256 425 2270
rect 375 2184 388 2256
rect 412 2184 425 2256
rect 375 2170 425 2184
rect 440 2256 490 2270
rect 440 2184 453 2256
rect 477 2184 490 2256
rect 440 2170 490 2184
rect 1876 2066 2076 2079
rect 1876 2045 1890 2066
rect 2057 2045 2076 2066
rect 1876 2029 2076 2045
rect -50 1983 0 2000
rect -50 16 -38 1983
rect -10 16 0 1983
rect -50 0 0 16
rect 2000 1980 2050 2000
rect 2000 13 2012 1980
rect 2040 13 2050 1980
rect 2000 0 2050 13
<< pdiff >>
rect 371 2608 971 2622
rect 371 2588 393 2608
rect 955 2588 971 2608
rect 371 2572 971 2588
rect -10 2485 290 2495
rect -10 2460 5 2485
rect 275 2460 290 2485
rect -10 2445 290 2460
rect 371 2528 971 2542
rect 371 2508 390 2528
rect 957 2508 971 2528
rect 371 2492 971 2508
rect -10 2233 290 2245
rect -10 2208 10 2233
rect 274 2208 290 2233
rect -10 2195 290 2208
rect 572 2194 1772 2204
rect 109 2140 159 2154
rect 109 2068 125 2140
rect 148 2068 159 2140
rect 109 2054 159 2068
rect 174 2141 224 2154
rect 174 2068 185 2141
rect 213 2068 224 2141
rect 572 2169 587 2194
rect 1757 2169 1772 2194
rect 572 2154 1772 2169
rect 174 2054 224 2068
rect 572 2092 1772 2104
rect 572 2067 587 2092
rect 1757 2067 1772 2092
rect 572 2054 1772 2067
<< ndiffc >>
rect 724 2403 1293 2428
rect 1395 2389 1807 2413
rect 1890 2393 2061 2419
rect 723 2323 1292 2348
rect 1395 2323 1807 2347
rect 388 2184 412 2256
rect 453 2184 477 2256
rect 1890 2045 2057 2066
rect -38 16 -10 1983
rect 2012 13 2040 1980
<< pdiffc >>
rect 393 2588 955 2608
rect 5 2460 275 2485
rect 390 2508 957 2528
rect 10 2208 274 2233
rect 125 2068 148 2140
rect 185 2068 213 2141
rect 587 2169 1757 2194
rect 587 2067 1757 2092
<< psubdiff >>
rect 2050 1985 2100 2000
rect 2050 15 2060 1985
rect 2090 15 2100 1985
rect 2050 0 2100 15
<< nsubdiff >>
rect 572 2234 1772 2255
rect 572 2213 587 2234
rect 1757 2213 1772 2234
rect 572 2204 1772 2213
rect 224 2141 274 2154
rect 224 2068 230 2141
rect 261 2068 274 2141
rect 224 2054 274 2068
<< psubdiffcont >>
rect 2060 15 2090 1985
<< nsubdiffcont >>
rect 587 2213 1757 2234
rect 230 2068 261 2141
<< poly >>
rect 358 2561 371 2572
rect 340 2542 371 2561
rect 971 2542 985 2572
rect 340 2468 355 2542
rect 340 2460 417 2468
rect 340 2453 389 2460
rect -23 2245 -10 2445
rect 290 2299 313 2445
rect 381 2436 389 2453
rect 409 2436 417 2460
rect 381 2428 417 2436
rect 687 2360 710 2390
rect 1310 2360 1324 2390
rect 1350 2375 1365 2437
rect 1350 2360 1375 2375
rect 1825 2360 1838 2375
rect 687 2299 702 2360
rect 290 2298 702 2299
rect 290 2283 712 2298
rect 290 2245 327 2283
rect 425 2282 712 2283
rect 425 2270 440 2282
rect 312 2177 327 2245
rect 159 2167 327 2177
rect 1861 2219 1876 2379
rect 159 2162 328 2167
rect 159 2154 174 2162
rect -40 2073 7 2083
rect -40 2043 -24 2073
rect -2 2043 7 2073
rect 295 2100 328 2162
rect 425 2157 440 2170
rect 1799 2211 1876 2219
rect 1799 2193 1808 2211
rect 1828 2193 1876 2211
rect 1799 2183 1876 2193
rect 551 2125 572 2154
rect 490 2105 572 2125
rect 390 2100 430 2105
rect 295 2095 430 2100
rect 295 2078 398 2095
rect 422 2078 430 2095
rect 295 2071 430 2078
rect 390 2069 430 2071
rect -40 2030 7 2043
rect 159 2038 174 2054
rect -40 2015 30 2030
rect 490 2015 508 2105
rect 551 2104 572 2105
rect 1772 2104 1785 2154
rect 1861 2104 1876 2183
rect 1860 2080 1876 2104
rect 1861 2079 1876 2080
rect 2076 2079 2100 2379
rect 1785 2058 1830 2070
rect 1785 2041 1796 2058
rect 1818 2041 1830 2058
rect 1785 2015 1830 2041
rect -40 2010 2000 2015
rect 0 2000 2000 2010
rect 0 -15 2000 0
<< polycont >>
rect 389 2436 409 2460
rect -24 2043 -2 2073
rect 1808 2193 1828 2211
rect 398 2078 422 2095
rect 1796 2041 1818 2058
<< locali >>
rect 1020 2615 1043 2619
rect 380 2608 1043 2615
rect 380 2588 393 2608
rect 955 2588 1043 2608
rect 380 2580 1043 2588
rect 1010 2557 1043 2580
rect 380 2528 965 2535
rect 380 2508 390 2528
rect 957 2508 965 2528
rect 380 2500 965 2508
rect -5 2485 285 2491
rect -5 2460 5 2485
rect 275 2460 285 2485
rect -5 2450 285 2460
rect 381 2460 416 2468
rect 381 2436 389 2460
rect 409 2436 416 2460
rect 595 2439 635 2500
rect 381 2265 416 2436
rect 594 2351 636 2439
rect 1010 2435 1044 2557
rect 715 2428 1305 2435
rect 715 2403 724 2428
rect 1293 2403 1305 2428
rect 1882 2419 2070 2423
rect 715 2395 1305 2403
rect 1385 2414 1815 2418
rect 1385 2389 1395 2414
rect 1807 2389 1815 2414
rect 1385 2382 1815 2389
rect 1882 2393 1890 2419
rect 2061 2393 2070 2419
rect 1882 2385 2070 2393
rect 715 2351 1305 2355
rect 594 2348 1305 2351
rect 594 2328 723 2348
rect 715 2323 723 2328
rect 1292 2323 1305 2348
rect 715 2315 1305 2323
rect 1385 2347 1815 2353
rect 1385 2323 1395 2347
rect 1807 2323 1815 2347
rect 1385 2317 1815 2323
rect 725 2298 765 2315
rect 380 2256 420 2265
rect -5 2233 285 2240
rect -5 2215 10 2233
rect -25 2208 10 2215
rect 274 2208 285 2233
rect 380 2214 388 2256
rect -25 2200 285 2208
rect -25 2083 7 2200
rect 340 2184 388 2214
rect 412 2184 420 2256
rect 340 2176 420 2184
rect -35 2073 7 2083
rect -35 2043 -24 2073
rect -2 2043 7 2073
rect -35 2033 7 2043
rect 119 2140 154 2149
rect 119 2068 125 2140
rect 148 2068 154 2140
rect 119 2059 154 2068
rect 179 2141 269 2149
rect 179 2068 185 2141
rect 213 2068 230 2141
rect 261 2068 269 2141
rect 179 2059 269 2068
rect 119 2040 150 2059
rect 340 2040 363 2176
rect 380 2175 420 2176
rect 445 2256 485 2265
rect 445 2184 453 2256
rect 477 2184 485 2256
rect 735 2244 775 2298
rect 1730 2244 1767 2317
rect 577 2234 1767 2244
rect 577 2213 587 2234
rect 1757 2213 1767 2234
rect 577 2201 1767 2213
rect 445 2175 485 2184
rect 578 2194 1767 2201
rect 578 2168 587 2194
rect 1757 2193 1767 2194
rect 1799 2211 1837 2219
rect 1799 2193 1808 2211
rect 1828 2193 1837 2211
rect 1757 2184 1837 2193
rect 1757 2169 1815 2184
rect 1757 2168 1767 2169
rect 578 2159 1767 2168
rect 390 2100 430 2105
rect 390 2099 580 2100
rect 390 2095 1767 2099
rect 390 2078 398 2095
rect 422 2092 1767 2095
rect 422 2082 587 2092
rect 422 2078 542 2082
rect 390 2072 542 2078
rect 390 2069 430 2072
rect 577 2067 587 2082
rect 1757 2067 1767 2092
rect 577 2059 1767 2067
rect 1785 2065 1830 2070
rect 1881 2066 2068 2075
rect 1881 2065 1890 2066
rect 119 2020 363 2040
rect 1785 2058 1890 2065
rect 1785 2041 1796 2058
rect 1818 2045 1890 2058
rect 2057 2045 2068 2066
rect 1818 2041 2068 2045
rect 1785 2035 2068 2041
rect 1785 2030 1830 2035
rect -45 1986 -5 1995
rect -45 16 -40 1986
rect -10 16 -5 1986
rect -45 5 -5 16
rect 2005 1985 2095 1995
rect 2005 1980 2060 1985
rect 2005 13 2012 1980
rect 2040 15 2060 1980
rect 2090 15 2095 1985
rect 2040 13 2095 15
rect 2005 5 2095 13
<< viali >>
rect 5 2460 275 2485
rect 1395 2413 1807 2414
rect 1395 2389 1807 2413
rect 1890 2393 2061 2419
rect 185 2068 211 2141
rect 230 2068 261 2141
rect 453 2184 477 2256
rect 587 2213 1757 2234
rect 587 2169 1757 2194
rect 587 2168 1757 2169
rect -40 1983 -10 1986
rect -40 16 -38 1983
rect -38 16 -10 1983
rect 2012 13 2040 1980
rect 2060 15 2090 1985
<< metal1 >>
rect 234 2639 989 2641
rect -10 2495 989 2639
rect -13 2485 989 2495
rect -13 2460 5 2485
rect 275 2481 989 2485
rect 275 2460 298 2481
rect -13 2446 298 2460
rect -13 2192 297 2446
rect 1375 2419 2091 2429
rect 1375 2414 1890 2419
rect 1375 2389 1395 2414
rect 1807 2393 1890 2414
rect 2061 2393 2091 2419
rect 1807 2389 2091 2393
rect 1375 2310 2091 2389
rect 1839 2284 2091 2310
rect 377 2270 424 2271
rect 374 2256 490 2270
rect -13 2190 281 2192
rect 107 2141 281 2190
rect 374 2184 453 2256
rect 477 2184 490 2256
rect 374 2169 490 2184
rect 571 2234 1772 2255
rect 571 2213 587 2234
rect 1757 2213 1772 2234
rect 571 2194 1772 2213
rect 107 2068 185 2141
rect 211 2068 230 2141
rect 261 2068 281 2141
rect 107 2048 281 2068
rect 377 2000 424 2169
rect 571 2168 587 2194
rect 1757 2168 1772 2194
rect 571 2054 1772 2168
rect 1840 2019 2091 2284
rect 1690 2000 2100 2019
rect -50 1986 2100 2000
rect -50 16 -40 1986
rect -10 1985 2100 1986
rect -10 1980 2060 1985
rect -10 16 2012 1980
rect -50 13 2012 16
rect 2040 15 2060 1980
rect 2090 15 2100 1985
rect 2040 13 2100 15
rect -50 -15 2100 13
<< labels >>
rlabel poly 1358 2437 1358 2437 1 W
port 1 n
rlabel poly 2100 2083 2100 2083 3 B
port 3 e
rlabel metal1 2100 2010 2100 2010 7 VN
port 2 w
rlabel poly -23 2304 -23 2304 7 A
port 4 w
rlabel metal1 -13 2484 -13 2484 7 VP
port 5 w
<< end >>
