magic
tech sky130A
magscale 1 2
timestamp 1702612896
<< nwell >>
rect -230 251 180 531
<< nmos >>
rect -120 -118 -90 82
rect 10 -118 40 82
rect 140 -118 170 82
rect 270 -118 300 82
<< pmos >>
rect 10 291 40 491
<< ndiff >>
rect -220 52 -120 82
rect -220 -88 -190 52
rect -150 -88 -120 52
rect -220 -118 -120 -88
rect -90 52 10 82
rect -90 -88 -60 52
rect -20 -88 10 52
rect -90 -118 10 -88
rect 40 52 140 82
rect 40 -88 70 52
rect 110 -88 140 52
rect 40 -118 140 -88
rect 170 52 270 82
rect 170 -88 200 52
rect 240 -88 270 52
rect 170 -118 270 -88
rect 300 52 400 82
rect 300 -88 330 52
rect 370 -88 400 52
rect 300 -118 400 -88
<< pdiff >>
rect -90 461 10 491
rect -90 321 -60 461
rect -20 321 10 461
rect -90 291 10 321
rect 40 461 140 491
rect 40 321 70 461
rect 110 321 140 461
rect 40 291 140 321
<< ndiffc >>
rect -190 -88 -150 52
rect -60 -88 -20 52
rect 70 -88 110 52
rect 200 -88 240 52
rect 330 -88 370 52
<< pdiffc >>
rect -60 321 -20 461
rect 70 321 110 461
<< psubdiff >>
rect -320 52 -220 82
rect -320 -88 -290 52
rect -250 -88 -220 52
rect -320 -118 -220 -88
rect 400 52 500 82
rect 400 -88 430 52
rect 470 -88 500 52
rect 400 -118 500 -88
<< nsubdiff >>
rect -190 461 -90 491
rect -190 321 -160 461
rect -120 321 -90 461
rect -190 291 -90 321
<< psubdiffcont >>
rect -290 -88 -250 52
rect 430 -88 470 52
<< nsubdiffcont >>
rect -160 321 -120 461
<< poly >>
rect 10 491 40 521
rect 170 301 250 321
rect 10 271 40 291
rect 170 271 190 301
rect 10 261 190 271
rect 230 261 250 301
rect 10 241 250 261
rect -40 172 40 192
rect -40 132 -20 172
rect 20 132 40 172
rect -40 112 170 132
rect -120 82 -90 112
rect 10 102 170 112
rect 10 82 40 102
rect 140 82 170 102
rect 270 82 300 112
rect -120 -148 -90 -118
rect -170 -168 -90 -148
rect -170 -208 -150 -168
rect -110 -208 -90 -168
rect -170 -228 -90 -208
rect 10 -148 40 -118
rect 140 -148 170 -118
rect 270 -148 300 -118
rect 10 -168 90 -148
rect 10 -208 30 -168
rect 70 -208 90 -168
rect 10 -228 90 -208
rect 270 -168 350 -148
rect 270 -208 290 -168
rect 330 -208 350 -168
rect 270 -228 350 -208
<< polycont >>
rect 190 261 230 301
rect -20 132 20 172
rect -150 -208 -110 -168
rect 30 -208 70 -168
rect 290 -208 330 -168
<< locali >>
rect -180 461 0 481
rect -180 321 -160 461
rect -120 321 -60 461
rect -20 321 0 461
rect -180 301 0 321
rect 50 461 130 481
rect 50 321 70 461
rect 110 341 130 461
rect 110 321 210 341
rect 50 301 250 321
rect 170 261 190 301
rect 230 261 250 301
rect 170 241 250 261
rect -40 172 40 192
rect -40 132 -20 172
rect 20 132 40 172
rect -40 112 40 132
rect -40 72 0 112
rect 180 72 220 241
rect -310 52 -130 72
rect -310 -88 -290 52
rect -250 -88 -190 52
rect -150 -88 -130 52
rect -310 -108 -130 -88
rect -80 52 0 72
rect -80 -88 -60 52
rect -20 -88 0 52
rect -80 -108 0 -88
rect 50 52 130 72
rect 50 -88 70 52
rect 110 -88 130 52
rect 50 -108 130 -88
rect 180 52 260 72
rect 180 -88 200 52
rect 240 -88 260 52
rect 180 -108 260 -88
rect 310 52 490 72
rect 310 -88 330 52
rect 370 -88 430 52
rect 470 -88 490 52
rect 310 -108 490 -88
rect -170 -148 -130 -108
rect 310 -148 350 -108
rect -170 -168 -90 -148
rect -170 -208 -150 -168
rect -110 -208 -90 -168
rect -170 -228 -90 -208
rect 10 -168 90 -148
rect 10 -208 30 -168
rect 70 -208 90 -168
rect 10 -228 90 -208
rect 270 -168 350 -148
rect 270 -208 290 -168
rect 330 -208 350 -168
rect 270 -228 350 -208
<< viali >>
rect -160 321 -120 461
rect -60 321 -20 461
rect -290 -88 -250 52
rect -190 -88 -150 52
rect 70 -88 110 52
rect 330 -88 370 52
rect 430 -88 470 52
<< metal1 >>
rect -190 461 140 491
rect -190 321 -160 461
rect -120 321 -60 461
rect -20 321 140 461
rect -190 291 140 321
rect -320 52 500 82
rect -320 -88 -290 52
rect -250 -88 -190 52
rect -150 -88 70 52
rect 110 -88 330 52
rect 370 -88 430 52
rect 470 -88 500 52
rect -320 -118 500 -88
<< labels >>
rlabel metal1 -190 391 -190 391 7 VP
port 1 w
rlabel locali 250 281 250 281 3 VBP
port 4 e
rlabel locali 50 -228 50 -228 5 VBN
port 3 s
rlabel metal1 -320 -18 -320 -18 7 VN
port 2 w
<< end >>
