magic
tech sky130A
timestamp 1702621683
<< poly >>
rect 2371 2444 2386 2449
rect 995 2285 1011 2322
rect 960 2262 1016 2285
rect 960 2136 975 2262
rect 925 2121 975 2136
rect 925 2090 945 2121
rect 3113 2115 3150 2116
rect 3113 2091 3155 2115
rect 890 2075 945 2090
rect 890 1794 905 2075
rect 865 1784 905 1794
rect 865 1764 875 1784
rect 895 1764 905 1784
rect 865 1754 905 1764
rect 3139 1522 3155 2091
rect 3139 1508 3265 1522
rect 3139 1504 3343 1508
rect 3139 1477 3366 1504
<< polycont >>
rect 875 1764 895 1784
<< locali >>
rect 865 1784 905 1794
rect 865 1764 875 1784
rect 895 1764 905 1784
rect 865 1754 905 1764
rect 4082 1753 4087 1772
rect 244 1479 248 1481
<< metal1 >>
rect 684 2649 789 2657
rect 1799 2650 3795 2654
rect 992 2649 3795 2650
rect 684 2646 3795 2649
rect 681 2634 3795 2646
rect 680 2548 3795 2634
rect 680 2029 789 2548
rect 992 2505 3795 2548
rect 992 2501 1828 2505
rect 41 1928 44 1934
rect 684 1829 789 2029
rect 3512 1947 3702 2505
rect 921 1734 925 1735
rect 880 1731 925 1734
rect 3115 1731 3216 1733
rect 41 1631 44 1637
rect 551 1536 3599 1731
rect 880 1534 925 1536
rect 921 1530 925 1534
rect 3115 1532 3216 1536
use memristor_emulator_res  memristor_emulator_res_0
timestamp 1702621296
transform 1 0 1021 0 1 12
box -100 -15 2100 2641
use neuron_top  neuron_top_0
timestamp 1702524960
transform 1 0 -28 0 1 1479
box -17 -1479 945 2073
use neuron_top  neuron_top_1
timestamp 1702524960
transform 1 0 3167 0 1 1477
box -17 -1479 945 2073
<< labels >>
rlabel metal1 42 1634 42 1634 3 VN
rlabel metal1 42 1929 42 1929 7 VP
rlabel poly 2379 2449 2379 2449 1 W
rlabel locali 4087 1763 4087 1763 3 VSYN
rlabel locali 247 1479 247 1479 5 ISYN
<< end >>
