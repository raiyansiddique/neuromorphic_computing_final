* NGSPICE file created from memristor_emulator_res.ext - technology: sky130A

.subckt memristor_emulator_res VP VN A B W
X0 VN B a_n80_4020# VN sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=3
X1 VN a_n80_4020# VN VN sky130_fd_pr__nfet_01v8 ad=10 pd=41 as=23.8 ps=100 w=20 l=20
X2 VP A a_n80_4020# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=2
X3 B a_n80_4020# A B sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=6 ps=25 w=12 l=0.5
X4 VP A a_218_4108# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X5 a_742_5144# A B VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.3
X6 a_742_5144# a_218_4108# B VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.3
X7 VN A a_218_4108# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X8 VN W B VN sky130_fd_pr__nfet_01v8 ad=2.25 pd=10 as=2.25 ps=10 w=4.5 l=0.15
.ends

