magic
tech sky130A
timestamp 1702324856
<< nwell >>
rect -48 2035 338 2371
rect 514 2160 1774 2400
<< nmos >>
rect 1876 2079 2076 2379
rect 0 0 2000 2000
<< pmos >>
rect 70 2053 270 2353
rect 544 2230 1744 2280
<< ndiff >>
rect 1876 2419 2076 2429
rect 1876 2393 1890 2419
rect 2061 2393 2076 2419
rect 1876 2379 2076 2393
rect 1876 2066 2076 2079
rect 1876 2045 1890 2066
rect 2057 2045 2076 2066
rect 1876 2029 2076 2045
rect -50 1983 0 2000
rect -50 16 -38 1983
rect -10 16 0 1983
rect -50 0 0 16
rect 2000 1980 2050 2000
rect 2000 13 2012 1980
rect 2040 13 2050 1980
rect 2000 0 2050 13
<< pdiff >>
rect 20 2338 70 2353
rect 20 2068 30 2338
rect 55 2068 70 2338
rect 20 2053 70 2068
rect 270 2337 320 2353
rect 270 2073 282 2337
rect 307 2073 320 2337
rect 544 2320 1744 2330
rect 544 2295 559 2320
rect 1729 2295 1744 2320
rect 544 2280 1744 2295
rect 270 2053 320 2073
rect 544 2218 1744 2230
rect 544 2193 559 2218
rect 1729 2193 1744 2218
rect 544 2180 1744 2193
<< ndiffc >>
rect 1890 2393 2061 2419
rect 1890 2045 2057 2066
rect -38 16 -10 1983
rect 2012 13 2040 1980
<< pdiffc >>
rect 30 2068 55 2338
rect 282 2073 307 2337
rect 559 2295 1729 2320
rect 559 2193 1729 2218
<< psubdiff >>
rect 2050 1985 2100 2000
rect 2050 15 2060 1985
rect 2090 15 2100 1985
rect 2050 0 2100 15
<< nsubdiff >>
rect -30 2338 20 2353
rect -30 2068 -15 2338
rect 10 2068 20 2338
rect -30 2053 20 2068
rect 544 2360 1744 2381
rect 544 2339 559 2360
rect 1729 2339 1744 2360
rect 544 2330 1744 2339
<< psubdiffcont >>
rect 2060 15 2090 1985
<< nsubdiffcont >>
rect -15 2068 10 2338
rect 559 2339 1729 2360
<< poly >>
rect 245 2376 386 2390
rect 70 2375 386 2376
rect 70 2353 270 2375
rect 369 2327 386 2375
rect 369 2324 410 2327
rect 370 2320 410 2324
rect 370 2303 378 2320
rect 401 2303 410 2320
rect 370 2295 410 2303
rect 1861 2327 1876 2379
rect 1799 2319 1876 2327
rect 1799 2301 1808 2319
rect 1828 2301 1876 2319
rect 1799 2291 1876 2301
rect 491 2230 544 2280
rect 1744 2230 1757 2280
rect 380 2171 430 2180
rect 380 2149 390 2171
rect 420 2149 430 2171
rect 70 2040 270 2053
rect 380 2015 430 2149
rect 490 2015 508 2230
rect 1861 2104 1876 2291
rect 1860 2080 1876 2104
rect 1861 2079 1876 2080
rect 2076 2079 2100 2379
rect 1785 2058 1830 2070
rect 1785 2041 1796 2058
rect 1818 2041 1830 2058
rect 1785 2015 1830 2041
rect 0 2000 2000 2015
rect 0 -15 2000 0
<< polycont >>
rect 378 2303 401 2320
rect 1808 2301 1828 2319
rect 390 2149 420 2171
rect 1796 2041 1818 2058
<< locali >>
rect 1882 2419 2070 2423
rect 1882 2393 1890 2419
rect 2061 2393 2070 2419
rect 1882 2385 2070 2393
rect 549 2360 1739 2370
rect -25 2338 65 2348
rect -25 2068 -15 2338
rect 10 2068 30 2338
rect 55 2068 65 2338
rect -25 2058 65 2068
rect 275 2337 315 2348
rect 275 2073 282 2337
rect 307 2180 315 2337
rect 549 2339 559 2360
rect 1729 2339 1739 2360
rect 549 2327 1739 2339
rect 370 2320 410 2327
rect 370 2303 378 2320
rect 401 2303 410 2320
rect 370 2295 410 2303
rect 390 2226 410 2295
rect 550 2320 1739 2327
rect 550 2294 559 2320
rect 1729 2319 1739 2320
rect 1799 2319 1837 2327
rect 1729 2301 1808 2319
rect 1828 2301 1837 2319
rect 1729 2295 1837 2301
rect 1729 2294 1739 2295
rect 550 2285 1739 2294
rect 1799 2292 1837 2295
rect 390 2225 552 2226
rect 390 2218 1739 2225
rect 390 2208 559 2218
rect 549 2193 559 2208
rect 1729 2193 1739 2218
rect 549 2185 1739 2193
rect 307 2171 430 2180
rect 307 2149 390 2171
rect 420 2149 430 2171
rect 307 2138 430 2149
rect 307 2073 315 2138
rect 275 2058 315 2073
rect 1785 2065 1830 2070
rect 1881 2066 2068 2075
rect 1881 2065 1890 2066
rect 1785 2058 1890 2065
rect 1785 2041 1796 2058
rect 1818 2045 1890 2058
rect 2057 2045 2068 2066
rect 1818 2041 2068 2045
rect 1785 2035 2068 2041
rect 1785 2030 1830 2035
rect -45 1986 -5 1995
rect -45 16 -40 1986
rect -10 16 -5 1986
rect -45 5 -5 16
rect 2005 1985 2095 1995
rect 2005 1980 2060 1985
rect 2005 13 2012 1980
rect 2040 15 2060 1980
rect 2090 15 2095 1985
rect 2040 13 2095 15
rect 2005 5 2095 13
<< viali >>
rect 1890 2393 2061 2419
rect -15 2068 10 2338
rect 30 2068 55 2338
rect 559 2339 1729 2360
rect 559 2295 1729 2320
rect 559 2294 1729 2295
rect -40 1983 -10 1986
rect -40 16 -38 1983
rect -38 16 -10 1983
rect 2012 13 2040 1980
rect 2060 15 2090 1985
<< metal1 >>
rect 1840 2419 2091 2429
rect 1840 2393 1890 2419
rect 2061 2393 2091 2419
rect 543 2360 1744 2381
rect -35 2338 325 2360
rect -35 2068 -15 2338
rect 10 2068 30 2338
rect 55 2068 325 2338
rect 543 2339 559 2360
rect 1729 2339 1744 2360
rect 543 2320 1744 2339
rect 543 2294 559 2320
rect 1729 2294 1744 2320
rect 543 2180 1744 2294
rect -35 2050 325 2068
rect 1840 2019 2091 2393
rect 1690 2000 2100 2019
rect -50 1986 2100 2000
rect -50 16 -40 1986
rect -10 1985 2100 1986
rect -10 1980 2060 1985
rect -10 16 2012 1980
rect -50 13 2012 16
rect 2040 15 2060 1980
rect 2090 15 2100 1985
rect 2040 13 2100 15
rect -50 -15 2100 13
<< labels >>
rlabel metal1 2100 2010 2100 2010 3 VN
rlabel poly 2100 2085 2100 2085 3 B
rlabel metal1 63 2360 63 2360 1 VP
rlabel poly 245 2385 245 2385 7 A
<< end >>
