magic
tech sky130A
timestamp 1702529013
<< poly >>
rect 2371 2444 2386 2449
rect 995 2285 1011 2322
rect 960 2262 1016 2285
rect 960 2136 975 2262
rect 925 2121 975 2136
rect 925 1794 942 2121
rect 3113 2115 3150 2116
rect 3113 2091 3155 2115
rect 910 1786 942 1794
rect 910 1762 917 1786
rect 936 1762 942 1786
rect 910 1754 942 1762
rect 3139 1522 3155 2091
rect 3139 1508 3265 1522
rect 3139 1504 3343 1508
rect 3139 1477 3366 1504
<< polycont >>
rect 917 1762 936 1786
<< locali >>
rect 891 1786 942 1794
rect 891 1762 917 1786
rect 936 1762 942 1786
rect 891 1754 942 1762
rect 4082 1753 4087 1772
rect 199 1479 203 1481
<< metal1 >>
rect 684 2649 789 2657
rect 1799 2650 3795 2654
rect 992 2649 3795 2650
rect 684 2646 3795 2649
rect 681 2634 3795 2646
rect 680 2548 3795 2634
rect 680 2029 789 2548
rect 992 2505 3795 2548
rect 992 2501 1828 2505
rect 41 1928 44 1934
rect 684 1829 789 2029
rect 3512 1947 3702 2505
rect 3115 1731 3216 1733
rect 41 1631 44 1637
rect 551 1536 3599 1731
rect 3115 1532 3216 1536
use memristor_emulator_res  memristor_emulator_res_0
timestamp 1702443510
transform 1 0 1021 0 1 12
box -50 -15 2100 2641
use neuron_top  neuron_top_0
timestamp 1702524960
transform 1 0 17 0 1 1479
box -17 -1479 945 2073
use neuron_top  neuron_top_1
timestamp 1702524960
transform 1 0 3167 0 1 1477
box -17 -1479 945 2073
<< labels >>
rlabel locali 4087 1763 4087 1763 3 VSYN
rlabel locali 202 1479 202 1479 5 ISYN
rlabel metal1 42 1634 42 1634 3 VN
rlabel metal1 42 1929 42 1929 7 VP
rlabel poly 2379 2449 2379 2449 1 W
<< end >>
