magic
tech sky130A
timestamp 1702431338
<< nwell >>
rect -48 2035 338 2371
rect 514 2050 1774 2290
<< nmos >>
rect 1876 2079 2076 2379
rect 0 0 2000 2000
<< pmos >>
rect 70 2053 270 2353
rect 544 2120 1744 2170
<< ndiff >>
rect 1876 2419 2076 2429
rect 1876 2393 1890 2419
rect 2061 2393 2076 2419
rect 1876 2379 2076 2393
rect 1876 2066 2076 2079
rect 1876 2045 1890 2066
rect 2057 2045 2076 2066
rect 1876 2029 2076 2045
rect -50 1983 0 2000
rect -50 16 -38 1983
rect -10 16 0 1983
rect -50 0 0 16
rect 2000 1980 2050 2000
rect 2000 13 2012 1980
rect 2040 13 2050 1980
rect 2000 0 2050 13
<< pdiff >>
rect 20 2338 70 2353
rect 20 2068 30 2338
rect 55 2068 70 2338
rect 20 2053 70 2068
rect 270 2337 320 2353
rect 270 2073 282 2337
rect 307 2073 320 2337
rect 544 2210 1744 2220
rect 544 2185 559 2210
rect 1729 2185 1744 2210
rect 270 2053 320 2073
rect 544 2170 1744 2185
rect 544 2108 1744 2120
rect 544 2083 559 2108
rect 1729 2083 1744 2108
rect 544 2070 1744 2083
<< ndiffc >>
rect 1890 2393 2061 2419
rect 1890 2045 2057 2066
rect -38 16 -10 1983
rect 2012 13 2040 1980
<< pdiffc >>
rect 30 2068 55 2338
rect 282 2073 307 2337
rect 559 2185 1729 2210
rect 559 2083 1729 2108
<< psubdiff >>
rect 2050 1985 2100 2000
rect 2050 15 2060 1985
rect 2090 15 2100 1985
rect 2050 0 2100 15
<< nsubdiff >>
rect -30 2338 20 2353
rect -30 2068 -15 2338
rect 10 2068 20 2338
rect -30 2053 20 2068
rect 544 2250 1744 2271
rect 544 2229 559 2250
rect 1729 2229 1744 2250
rect 544 2220 1744 2229
<< psubdiffcont >>
rect 2060 15 2090 1985
<< nsubdiffcont >>
rect -15 2068 10 2338
rect 559 2229 1729 2250
<< poly >>
rect 245 2376 386 2390
rect 70 2375 386 2376
rect 70 2353 270 2375
rect 369 2327 386 2375
rect 369 2324 410 2327
rect 370 2320 410 2324
rect 370 2303 378 2320
rect 401 2303 410 2320
rect 370 2295 410 2303
rect 1861 2219 1876 2379
rect 380 2171 430 2180
rect 380 2149 390 2171
rect 420 2149 430 2171
rect 1799 2211 1876 2219
rect 1799 2193 1808 2211
rect 1828 2193 1876 2211
rect 1799 2183 1876 2193
rect 70 2040 270 2053
rect 380 2015 430 2149
rect 491 2120 544 2170
rect 1744 2120 1757 2170
rect 490 2015 508 2120
rect 1861 2104 1876 2183
rect 1860 2080 1876 2104
rect 1861 2079 1876 2080
rect 2076 2079 2100 2379
rect 1785 2058 1830 2070
rect 1785 2041 1796 2058
rect 1818 2041 1830 2058
rect 1785 2015 1830 2041
rect 0 2000 2000 2015
rect 0 -15 2000 0
<< polycont >>
rect 378 2303 401 2320
rect 390 2149 420 2171
rect 1808 2193 1828 2211
rect 1796 2041 1818 2058
<< locali >>
rect 1882 2419 2070 2423
rect 1882 2393 1890 2419
rect 2061 2393 2070 2419
rect 1882 2385 2070 2393
rect -25 2338 65 2348
rect -25 2068 -15 2338
rect 10 2068 30 2338
rect 55 2068 65 2338
rect -25 2058 65 2068
rect 275 2337 315 2348
rect 275 2073 282 2337
rect 307 2180 315 2337
rect 370 2320 410 2327
rect 370 2303 378 2320
rect 401 2303 410 2320
rect 370 2295 410 2303
rect 390 2226 410 2295
rect 549 2250 1739 2260
rect 549 2229 559 2250
rect 1729 2229 1739 2250
rect 477 2226 495 2229
rect 390 2208 495 2226
rect 549 2217 1739 2229
rect 307 2171 430 2180
rect 307 2149 390 2171
rect 420 2149 430 2171
rect 307 2138 430 2149
rect 307 2073 315 2138
rect 477 2116 495 2208
rect 550 2210 1739 2217
rect 1799 2211 1837 2219
rect 550 2184 559 2210
rect 1729 2209 1739 2210
rect 1793 2209 1808 2211
rect 1729 2193 1808 2209
rect 1828 2193 1837 2211
rect 1729 2185 1837 2193
rect 1729 2184 1739 2185
rect 1771 2184 1837 2185
rect 550 2175 1739 2184
rect 477 2115 552 2116
rect 477 2108 1739 2115
rect 477 2099 559 2108
rect 478 2098 559 2099
rect 549 2083 559 2098
rect 1729 2083 1739 2108
rect 549 2075 1739 2083
rect 275 2058 315 2073
rect 1785 2065 1830 2070
rect 1881 2066 2068 2075
rect 1881 2065 1890 2066
rect 1785 2058 1890 2065
rect 1785 2041 1796 2058
rect 1818 2045 1890 2058
rect 2057 2045 2068 2066
rect 1818 2041 2068 2045
rect 1785 2035 2068 2041
rect 1785 2030 1830 2035
rect -45 1986 -5 1995
rect -45 16 -40 1986
rect -10 16 -5 1986
rect -45 5 -5 16
rect 2005 1985 2095 1995
rect 2005 1980 2060 1985
rect 2005 13 2012 1980
rect 2040 15 2060 1980
rect 2090 15 2095 1985
rect 2040 13 2095 15
rect 2005 5 2095 13
<< viali >>
rect 1890 2393 2061 2419
rect -15 2068 10 2338
rect 30 2068 55 2338
rect 559 2229 1729 2250
rect 559 2185 1729 2210
rect 559 2184 1729 2185
rect -40 1983 -10 1986
rect -40 16 -38 1983
rect -38 16 -10 1983
rect 2012 13 2040 1980
rect 2060 15 2090 1985
<< metal1 >>
rect 1840 2419 2091 2429
rect 1840 2393 1890 2419
rect 2061 2393 2091 2419
rect -35 2338 325 2360
rect -35 2068 -15 2338
rect 10 2068 30 2338
rect 55 2068 325 2338
rect 1840 2331 2091 2393
rect 1861 2291 2091 2331
rect 543 2250 1744 2271
rect 543 2229 559 2250
rect 1729 2229 1744 2250
rect 543 2210 1744 2229
rect 543 2184 559 2210
rect 1729 2184 1744 2210
rect 543 2070 1744 2184
rect -35 2050 325 2068
rect 1840 2019 2091 2291
rect 1690 2000 2100 2019
rect -50 1986 2100 2000
rect -50 16 -40 1986
rect -10 1985 2100 1986
rect -10 1980 2060 1985
rect -10 16 2012 1980
rect -50 13 2012 16
rect 2040 15 2060 1980
rect 2090 15 2100 1985
rect 2040 13 2100 15
rect -50 -15 2100 13
<< labels >>
rlabel metal1 2100 2010 2100 2010 3 VN
port 3 e
rlabel poly 2100 2085 2100 2085 3 B
port 2 e
rlabel metal1 63 2360 63 2360 1 VP
port 4 n
rlabel poly 245 2385 245 2385 7 A
port 1 w
<< end >>
