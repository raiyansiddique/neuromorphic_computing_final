magic
tech sky130A
timestamp 1702075234
<< nwell >>
rect -95 -25 765 215
<< nmos >>
rect -25 -300 5 -100
rect 55 -300 85 -100
rect 215 -300 245 -100
rect 295 -300 325 -100
rect 455 -300 485 -100
rect 535 -300 565 -100
rect 745 -300 775 -100
<< pmos >>
rect -25 -5 5 195
rect 55 -5 85 195
rect 135 -5 165 195
rect 215 -5 245 195
rect 375 -5 405 195
rect 455 -5 485 195
rect 665 -5 695 195
<< ndiff >>
rect -75 -115 -25 -100
rect -75 -285 -60 -115
rect -40 -285 -25 -115
rect -75 -300 -25 -285
rect 5 -115 55 -100
rect 5 -285 20 -115
rect 40 -285 55 -115
rect 5 -300 55 -285
rect 85 -115 135 -100
rect 85 -285 100 -115
rect 120 -285 135 -115
rect 85 -300 135 -285
rect 165 -115 215 -100
rect 165 -285 180 -115
rect 200 -285 215 -115
rect 165 -300 215 -285
rect 245 -115 295 -100
rect 245 -285 260 -115
rect 280 -285 295 -115
rect 245 -300 295 -285
rect 325 -115 375 -100
rect 325 -285 340 -115
rect 360 -285 375 -115
rect 325 -300 375 -285
rect 405 -115 455 -100
rect 405 -285 420 -115
rect 440 -285 455 -115
rect 405 -300 455 -285
rect 485 -115 535 -100
rect 485 -285 500 -115
rect 520 -285 535 -115
rect 485 -300 535 -285
rect 565 -115 615 -100
rect 565 -285 580 -115
rect 600 -285 615 -115
rect 565 -300 615 -285
rect 695 -115 745 -100
rect 695 -285 710 -115
rect 730 -285 745 -115
rect 695 -300 745 -285
rect 775 -115 825 -100
rect 775 -285 790 -115
rect 810 -285 825 -115
rect 775 -300 825 -285
<< pdiff >>
rect -75 180 -25 195
rect -75 10 -60 180
rect -40 10 -25 180
rect -75 -5 -25 10
rect 5 180 55 195
rect 5 10 20 180
rect 40 10 55 180
rect 5 -5 55 10
rect 85 180 135 195
rect 85 10 100 180
rect 120 10 135 180
rect 85 -5 135 10
rect 165 180 215 195
rect 165 10 180 180
rect 200 10 215 180
rect 165 -5 215 10
rect 245 180 295 195
rect 245 10 260 180
rect 280 10 295 180
rect 245 -5 295 10
rect 325 180 375 195
rect 325 10 340 180
rect 360 10 375 180
rect 325 -5 375 10
rect 405 180 455 195
rect 405 10 420 180
rect 440 10 455 180
rect 405 -5 455 10
rect 485 180 535 195
rect 485 10 500 180
rect 520 10 535 180
rect 485 -5 535 10
rect 615 180 665 195
rect 615 10 630 180
rect 650 10 665 180
rect 615 -5 665 10
rect 695 180 745 195
rect 695 10 710 180
rect 730 10 745 180
rect 695 -5 745 10
<< ndiffc >>
rect -60 -285 -40 -115
rect 20 -285 40 -115
rect 100 -285 120 -115
rect 180 -285 200 -115
rect 260 -285 280 -115
rect 340 -285 360 -115
rect 420 -285 440 -115
rect 500 -285 520 -115
rect 580 -285 600 -115
rect 710 -285 730 -115
rect 790 -285 810 -115
<< pdiffc >>
rect -60 10 -40 180
rect 20 10 40 180
rect 100 10 120 180
rect 180 10 200 180
rect 260 10 280 180
rect 340 10 360 180
rect 420 10 440 180
rect 500 10 520 180
rect 630 10 650 180
rect 710 10 730 180
<< psubdiff >>
rect 645 -115 695 -100
rect 645 -285 660 -115
rect 680 -285 695 -115
rect 645 -300 695 -285
<< nsubdiff >>
rect 565 180 615 195
rect 565 10 580 180
rect 600 10 615 180
rect 565 -5 615 10
<< psubdiffcont >>
rect 660 -285 680 -115
<< nsubdiffcont >>
rect 580 10 600 180
<< poly >>
rect 135 240 175 250
rect 135 220 145 240
rect 165 220 175 240
rect 135 210 175 220
rect 365 240 405 250
rect 365 220 375 240
rect 395 220 405 240
rect 365 210 405 220
rect -25 195 5 210
rect 55 195 85 210
rect 135 195 165 210
rect 215 195 245 210
rect 375 195 405 210
rect 455 195 485 210
rect 665 195 695 210
rect -25 -15 5 -5
rect 55 -15 85 -5
rect -25 -20 85 -15
rect 135 -20 165 -5
rect 215 -20 245 -5
rect 375 -20 405 -5
rect 455 -20 485 -5
rect 665 -20 695 -5
rect -50 -30 85 -20
rect 205 -30 245 -20
rect -50 -50 -40 -30
rect -20 -50 -10 -30
rect -50 -60 -10 -50
rect 205 -50 215 -30
rect 235 -45 245 -30
rect 390 -35 430 -20
rect 235 -50 310 -45
rect 205 -60 310 -50
rect 295 -85 310 -60
rect 415 -75 430 -35
rect 470 -35 485 -20
rect 470 -50 550 -35
rect 415 -85 470 -75
rect 535 -85 550 -50
rect 610 -55 650 -45
rect 610 -75 620 -55
rect 640 -70 650 -55
rect 680 -70 695 -20
rect 640 -75 760 -70
rect 610 -85 760 -75
rect -25 -100 5 -85
rect 55 -100 85 -85
rect 215 -100 245 -85
rect 295 -100 325 -85
rect 415 -90 485 -85
rect 455 -100 485 -90
rect 535 -100 565 -85
rect 745 -100 775 -85
rect -25 -310 5 -300
rect 55 -310 85 -300
rect -25 -315 85 -310
rect 215 -315 245 -300
rect 295 -315 325 -300
rect 455 -315 485 -300
rect 535 -315 565 -300
rect 745 -315 775 -300
rect -25 -325 110 -315
rect 70 -345 80 -325
rect 100 -345 110 -325
rect 70 -355 110 -345
rect 215 -325 255 -315
rect 215 -345 225 -325
rect 245 -345 255 -325
rect 215 -355 255 -345
rect 525 -325 565 -315
rect 525 -345 535 -325
rect 555 -345 565 -325
rect 525 -355 565 -345
<< polycont >>
rect 145 220 165 240
rect 375 220 395 240
rect -40 -50 -20 -30
rect 215 -50 235 -30
rect 620 -75 640 -55
rect 80 -345 100 -325
rect 225 -345 245 -325
rect 535 -345 555 -325
<< locali >>
rect 135 240 175 250
rect 135 220 145 240
rect 165 230 175 240
rect 365 240 405 250
rect 365 230 375 240
rect 165 220 375 230
rect 395 220 405 240
rect 135 210 405 220
rect 250 190 270 210
rect -70 180 -30 190
rect -70 10 -60 180
rect -40 10 -30 180
rect -70 0 -30 10
rect 10 180 50 190
rect 10 10 20 180
rect 40 10 50 180
rect 10 0 50 10
rect 90 180 130 190
rect 90 10 100 180
rect 120 10 130 180
rect 90 0 130 10
rect 170 180 210 190
rect 170 10 180 180
rect 200 10 210 180
rect 170 0 210 10
rect 250 180 290 190
rect 250 10 260 180
rect 280 10 290 180
rect 250 0 290 10
rect -50 -20 -30 0
rect 110 -20 130 0
rect -50 -30 -10 -20
rect -50 -50 -40 -30
rect -20 -50 -10 -30
rect 110 -30 245 -20
rect 110 -40 215 -30
rect -50 -60 -10 -50
rect 190 -50 215 -40
rect 235 -50 245 -30
rect 190 -60 245 -50
rect 270 -60 290 0
rect 330 180 370 190
rect 330 10 340 180
rect 360 10 370 180
rect 330 0 370 10
rect 410 180 450 190
rect 410 10 420 180
rect 440 10 450 180
rect 410 0 450 10
rect 490 180 530 190
rect 490 10 500 180
rect 520 10 530 180
rect 490 0 530 10
rect 570 180 660 190
rect 570 10 580 180
rect 600 10 630 180
rect 650 10 660 180
rect 570 0 660 10
rect 700 180 740 190
rect 700 10 710 180
rect 730 10 740 180
rect 700 0 740 10
rect 330 -20 350 0
rect 510 -20 530 0
rect 330 -40 410 -20
rect 510 -40 590 -20
rect -50 -105 -30 -60
rect 190 -105 210 -60
rect 270 -80 350 -60
rect 330 -105 350 -80
rect 390 -80 410 -40
rect 570 -45 590 -40
rect 720 -40 740 0
rect 570 -55 650 -45
rect 570 -65 620 -55
rect 390 -100 430 -80
rect 410 -105 430 -100
rect 570 -105 590 -65
rect 610 -75 620 -65
rect 640 -75 650 -55
rect 720 -60 800 -40
rect 610 -85 650 -75
rect 780 -80 825 -60
rect 780 -105 800 -80
rect -70 -115 -30 -105
rect -70 -285 -60 -115
rect -40 -285 -30 -115
rect -70 -295 -30 -285
rect 10 -115 50 -105
rect 10 -285 20 -115
rect 40 -285 50 -115
rect 10 -295 50 -285
rect 90 -115 130 -105
rect 90 -285 100 -115
rect 120 -285 130 -115
rect 90 -295 130 -285
rect 170 -115 210 -105
rect 170 -285 180 -115
rect 200 -285 210 -115
rect 170 -295 210 -285
rect 250 -115 290 -105
rect 250 -285 260 -115
rect 280 -285 290 -115
rect 250 -295 290 -285
rect 330 -115 370 -105
rect 330 -285 340 -115
rect 360 -285 370 -115
rect 330 -295 370 -285
rect 410 -115 450 -105
rect 410 -285 420 -115
rect 440 -285 450 -115
rect 410 -295 450 -285
rect 490 -115 530 -105
rect 490 -285 500 -115
rect 520 -285 530 -115
rect 490 -295 530 -285
rect 570 -115 610 -105
rect 570 -285 580 -115
rect 600 -285 610 -115
rect 570 -295 610 -285
rect 650 -115 740 -105
rect 650 -285 660 -115
rect 680 -285 710 -115
rect 730 -285 740 -115
rect 650 -295 740 -285
rect 780 -115 820 -105
rect 780 -285 790 -115
rect 810 -285 820 -115
rect 780 -295 820 -285
rect 90 -315 110 -295
rect 410 -315 430 -295
rect 70 -325 110 -315
rect 70 -345 80 -325
rect 100 -345 110 -325
rect 70 -355 110 -345
rect 215 -325 565 -315
rect 215 -345 225 -325
rect 245 -335 535 -325
rect 245 -345 255 -335
rect 215 -355 255 -345
rect 525 -345 535 -335
rect 555 -345 565 -325
rect 525 -355 565 -345
<< viali >>
rect 20 10 40 180
rect 180 10 200 180
rect 420 10 440 180
rect 580 10 600 180
rect 630 10 650 180
rect 20 -285 40 -115
rect 260 -285 280 -115
rect 500 -285 520 -115
rect 660 -285 680 -115
rect 710 -285 730 -115
<< metal1 >>
rect -75 180 745 195
rect -75 10 20 180
rect 40 10 180 180
rect 200 10 420 180
rect 440 10 580 180
rect 600 10 630 180
rect 650 10 745 180
rect -75 -5 745 10
rect -75 -115 825 -100
rect -75 -285 20 -115
rect 40 -285 260 -115
rect 280 -285 500 -115
rect 520 -285 660 -115
rect 680 -285 710 -115
rect 730 -285 825 -115
rect -75 -300 825 -285
<< labels >>
rlabel metal1 -70 95 -70 95 7 VP
rlabel metal1 -70 -200 -70 -200 7 VN
rlabel locali 90 -355 90 -355 5 IEX
rlabel locali 825 -70 825 -70 3 VOUT
<< end >>
